-- Memory (512 x 16)

library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.STD_LOGIC_UNSIGNED.ALL;

entity memory is
	port(
		data_I, addr_I: in std_logic_vector (15 downto 0);
		MW: in std_logic;
		data_O: out std_logic_vector (15 downto 0)
	);
end memory;

architecture behave of memory is
	type mem_array is array(0 to 511) of std_logic_vector (15 downto 0);
begin
	mem_process: process(addr_I, data_I, MW)
	variable mem: mem_array := (
		-- 00
		x"1337", x"DEAD", x"BEEF", x"000F",
		x"0000", x"0000", x"0000", x"0000",
		x"0000", x"0000", x"0000", x"0000",
		x"0000", x"0000", x"0000", x"0000",
		-- 01
		x"0000", x"0000", x"0000", x"0000",
		x"0000", x"0000", x"0000", x"0000",
		x"0000", x"0000", x"0000", x"0000",
		x"0000", x"0000", x"0000", x"0000",
		-- 02
		x"0000", x"0000", x"0000", x"0000",
		x"0000", x"0000", x"0000", x"0000",
		x"0000", x"0000", x"0000", x"0000",
		x"0000", x"0000", x"0000", x"0000",
		-- 03
		x"0000", x"0000", x"0000", x"0000",
		x"0000", x"0000", x"0000", x"0000",
		x"0000", x"0000", x"0000", x"0000",
		x"0000", x"0000", x"0000", x"0000",
		-- 04
		x"0000", x"0000", x"0000", x"0000",
		x"0000", x"0000", x"0000", x"0000",
		x"0000", x"0000", x"0000", x"0000",
		x"0000", x"0000", x"0000", x"0000",
		-- 05
		x"0000", x"0000", x"0000", x"0000",
		x"0000", x"0000", x"0000", x"0000",
		x"0000", x"0000", x"0000", x"0000",
		x"0000", x"0000", x"0000", x"0000",
		-- 06
		x"0000", x"0000", x"0000", x"0000",
		x"0000", x"0000", x"0000", x"0000",
		x"0000", x"0000", x"0000", x"0000",
		x"0000", x"0000", x"0000", x"0000",
		-- 07
		x"0000", x"0000", x"0000", x"0000",
		x"0000", x"0000", x"0000", x"0000",
		x"0000", x"0000", x"0000", x"0000",
		x"0000", x"0000", x"0000", x"0000",
		-- 08
		x"0000", x"0000", x"0000", x"0000",
		x"0000", x"0000", x"0000", x"0000",
		x"0000", x"0000", x"0000", x"0000",
		x"0000", x"0000", x"0000", x"0000",
		-- 09
		x"0000", x"0000", x"0000", x"0000",
		x"0000", x"0000", x"0000", x"0000",
		x"0000", x"0000", x"0000", x"0000",
		x"0000", x"0000", x"0000", x"0000",
		-- 0A
		x"0000", x"0000", x"0000", x"0000",
		x"0000", x"0000", x"0000", x"0000",
		x"0000", x"0000", x"0000", x"0000",
		x"0000", x"0000", x"0000", x"0000",
		-- 0B
		x"0000", x"0000", x"0000", x"0000",
		x"0000", x"0000", x"0000", x"0000",
		x"0000", x"0000", x"0000", x"0000",
		x"0000", x"0000", x"0000", x"0000",
		-- 0C
		x"0000", x"0000", x"0000", x"0000",
		x"0000", x"0000", x"0000", x"0000",
		x"0000", x"0000", x"0000", x"0000",
		x"0000", x"0000", x"0000", x"0000",
		-- 0D
		x"0000", x"0000", x"0000", x"0000",
		x"0000", x"0000", x"0000", x"0000",
		x"0000", x"0000", x"0000", x"0000",
		x"0000", x"0000", x"0000", x"0000",
		-- 0E
		x"0000", x"0000", x"0000", x"0000",
		x"0000", x"0000", x"0000", x"0000",
		x"0000", x"0000", x"0000", x"0000",
		x"0000", x"0000", x"0000", x"0000",
		-- 0F
		x"0000", x"0000", x"0000", x"0000",
		x"0000", x"0000", x"0000", x"0000",
		x"0000", x"0000", x"0000", x"0000",
		x"0000", x"0000", x"0000", x"0000",
		-- 10
		x"0000", x"0000", x"0000", x"0000",
		x"0000", x"0000", x"0000", x"0000",
		x"0000", x"0000", x"0000", x"0000",
		x"0000", x"0000", x"0000", x"0000",
		-- 11
		x"0000", x"0000", x"0000", x"0000",
		x"0000", x"0000", x"0000", x"0000",
		x"0000", x"0000", x"0000", x"0000",
		x"0000", x"0000", x"0000", x"0000",
		-- 12
		x"0000", x"0000", x"0000", x"0000",
		x"0000", x"0000", x"0000", x"0000",
		x"0000", x"0000", x"0000", x"0000",
		x"0000", x"0000", x"0000", x"0000",
		-- 13
		x"0000", x"0000", x"0000", x"0000",
		x"0000", x"0000", x"0000", x"0000",
		x"0000", x"0000", x"0000", x"0000",
		x"0000", x"0000", x"0000", x"0000",
		-- 14
		x"0000", x"0000", x"0000", x"0000",
		x"0000", x"0000", x"0000", x"0000",
		x"0000", x"0000", x"0000", x"0000",
		x"0000", x"0000", x"0000", x"0000",
		-- 15
		x"0000", x"0000", x"0000", x"0000",
		x"0000", x"0000", x"0000", x"0000",
		x"0000", x"0000", x"0000", x"0000",
		x"0000", x"0000", x"0000", x"0000",
		-- 16
		x"0000", x"0000", x"0000", x"0000",
		x"0000", x"0000", x"0000", x"0000",
		x"0000", x"0000", x"0000", x"0000",
		x"0000", x"0000", x"0000", x"0000",
		-- 17
		x"0000", x"0000", x"0000", x"0000",
		x"0000", x"0000", x"0000", x"0000",
		x"0000", x"0000", x"0000", x"0000",
		x"0000", x"0000", x"0000", x"0000",
		-- 18
		x"0000", x"0000", x"0000", x"0000",
		x"0000", x"0000", x"0000", x"0000",
		x"0000", x"0000", x"0000", x"0000",
		x"0000", x"0000", x"0000", x"0000",
		-- 19
		x"0000", x"0000", x"0000", x"0000",
		x"0000", x"0000", x"0000", x"0000",
		x"0000", x"0000", x"0000", x"0000",
		x"0000", x"0000", x"0000", x"0000",
		-- 1A
		x"0000", x"0000", x"0000", x"0000",
		x"0000", x"0000", x"0000", x"0000",
		x"0000", x"0000", x"0000", x"0000",
		x"0000", x"0000", x"0000", x"0000",
		-- 1B
		x"0000", x"0000", x"0000", x"0000",
		x"0000", x"0000", x"0000", x"0000",
		x"0000", x"0000", x"0000", x"0000",
		x"0000", x"0000", x"0000", x"0000",
		-- 1C
		x"0000", x"0000", x"0000", x"0000",
		x"0000", x"0000", x"0000", x"0000",
		x"0000", x"0000", x"0000", x"0000",
		x"0000", x"0000", x"0000", x"0000",
		-- 1D
		x"0000", x"0000", x"0000", x"0000",
		x"0000", x"0000", x"0000", x"0000",
		x"0000", x"0000", x"0000", x"0000",
		x"0000", x"0000", x"0000", x"0000",
		-- 1E
		x"0000", x"0000", x"0000", x"0000",
		x"0000", x"0000", x"0000", x"0000",
		x"0000", x"0000", x"0000", x"0000",
		x"0000", x"0000", x"0000", x"0000",
		-- 1F
		x"0000", x"0000", x"0000", x"0000",
		x"0000", x"0000", x"0000", x"0000",
		x"0000", x"0000", x"0000", x"0000",
		x"0000", x"0000", x"0000", x"0000"
	);

	variable addr_C: integer range 0 to 511;
	variable addr_O: std_logic_vector(15 downto 0);

	begin
		
		addr_C := conv_integer(addr_I(8 downto 0));
		addr_O := mem(addr_C);
		
		if MW = '1' then mem(addr_C) := data_I;
		else data_O <= addr_O;
		end if;

	end process;
	
end behave;
