-- Datapath (TLS)

library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
